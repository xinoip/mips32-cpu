`define DELAY 20
module equal_32_testbench();
	reg [31:0] a, b;
    wire result;
	
    equal_32 test_equal_32(result, a, b);
	
initial begin
	a = 32'b00000000000000000000000000000000;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b11111111111111111111111111111111;
    b = 32'b11111111111111111111111111111111;
#`DELAY;
    a = 32'b00000000000000000000000000000001;
    b = 32'b00000000000000000000000000000000;
#`DELAY;
    a = 32'b00000000000001000000000000000000;
    b = 32'b00000000010000010000000000000000;
#`DELAY;
    a = 32'b10000000010001010001110000000000;
    b = 32'b10000000010001010001110000000000;
#`DELAY;
end

initial begin
	$monitor("time=%2d, a=%32b, b=%32b, result=%1b", $time, a, b, result);
end

endmodule
	