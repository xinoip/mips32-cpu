module mux32x4 (result, i0, i1, i2, i3, select);
    input [31:0] i0, i1, i2, i3;
    input [1:0] select;
    output [31:0] result;

    mux4 m1(result[0], i0[0], i1[0], i2[0], i3[0], select);
    mux4 m2(result[1], i0[1], i1[1], i2[1], i3[1], select);
    mux4 m3(result[2], i0[2], i1[2], i2[2], i3[2], select);
    mux4 m4(result[3], i0[3], i1[3], i2[3], i3[3], select);
    mux4 m5(result[4], i0[4], i1[4], i2[4], i3[4], select);
    mux4 m6(result[5], i0[5], i1[5], i2[5], i3[5], select);
    mux4 m7(result[6], i0[6], i1[6], i2[6], i3[6], select);
    mux4 m8(result[7], i0[7], i1[7], i2[7], i3[7], select);
    mux4 m9(result[8], i0[8], i1[8], i2[8], i3[8], select);
    mux4 m10(result[9], i0[9], i1[9], i2[9], i3[9], select);
    mux4 m11(result[10], i0[10], i1[10], i2[10], i3[10], select);
    mux4 m12(result[11], i0[11], i1[11], i2[11], i3[11], select);
    mux4 m13(result[12], i0[12], i1[12], i2[12], i3[12], select);
    mux4 m14(result[13], i0[13], i1[13], i2[13], i3[13], select);
    mux4 m15(result[14], i0[14], i1[14], i2[14], i3[14], select);
    mux4 m16(result[15], i0[15], i1[15], i2[15], i3[15], select);
    mux4 m17(result[16], i0[16], i1[16], i2[16], i3[16], select);
    mux4 m18(result[17], i0[17], i1[17], i2[17], i3[17], select);
    mux4 m19(result[18], i0[18], i1[18], i2[18], i3[18], select);
    mux4 m20(result[19], i0[19], i1[19], i2[19], i3[19], select);
    mux4 m21(result[20], i0[20], i1[20], i2[20], i3[20], select);
    mux4 m22(result[21], i0[21], i1[21], i2[21], i3[21], select);
    mux4 m23(result[22], i0[22], i1[22], i2[22], i3[22], select);
    mux4 m24(result[23], i0[23], i1[23], i2[23], i3[23], select);
    mux4 m25(result[24], i0[24], i1[24], i2[24], i3[24], select);
    mux4 m26(result[25], i0[25], i1[25], i2[25], i3[25], select);
    mux4 m27(result[26], i0[26], i1[26], i2[26], i3[26], select);
    mux4 m28(result[27], i0[27], i1[27], i2[27], i3[27], select);
    mux4 m29(result[28], i0[28], i1[28], i2[28], i3[28], select);
    mux4 m30(result[29], i0[29], i1[29], i2[29], i3[29], select);
    mux4 m31(result[30], i0[30], i1[30], i2[30], i3[30], select);
    mux4 m32(result[31], i0[31], i1[31], i2[31], i3[31], select);
endmodule