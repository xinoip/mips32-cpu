module mux32x2 (result, i0, i1, select);
    input [31:0] i0, i1;
    output [31:0] result;
    input select;

    mux2 m1(result[0], i0[0], i1[0], select);
    mux2 m2(result[1], i0[1], i1[1], select);
    mux2 m3(result[2], i0[2], i1[2], select);
    mux2 m4(result[3], i0[3], i1[3], select);
    mux2 m5(result[4], i0[4], i1[4], select);
    mux2 m6(result[5], i0[5], i1[5], select);
    mux2 m7(result[6], i0[6], i1[6], select);
    mux2 m8(result[7], i0[7], i1[7], select);
    mux2 m9(result[8], i0[8], i1[8], select);
    mux2 m10(result[9], i0[9], i1[9], select);
    mux2 m11(result[10], i0[10], i1[10], select);
    mux2 m12(result[11], i0[11], i1[11], select);
    mux2 m13(result[12], i0[12], i1[12], select);
    mux2 m14(result[13], i0[13], i1[13], select);
    mux2 m15(result[14], i0[14], i1[14], select);
    mux2 m16(result[15], i0[15], i1[15], select);
    mux2 m17(result[16], i0[16], i1[16], select);
    mux2 m18(result[17], i0[17], i1[17], select);
    mux2 m19(result[18], i0[18], i1[18], select);
    mux2 m20(result[19], i0[19], i1[19], select);
    mux2 m21(result[20], i0[20], i1[20], select);
    mux2 m22(result[21], i0[21], i1[21], select);
    mux2 m23(result[22], i0[22], i1[22], select);
    mux2 m24(result[23], i0[23], i1[23], select);
    mux2 m25(result[24], i0[24], i1[24], select);
    mux2 m26(result[25], i0[25], i1[25], select);
    mux2 m27(result[26], i0[26], i1[26], select);
    mux2 m28(result[27], i0[27], i1[27], select);
    mux2 m29(result[28], i0[28], i1[28], select);
    mux2 m30(result[29], i0[29], i1[29], select);
    mux2 m31(result[30], i0[30], i1[30], select);
    mux2 m32(result[31], i0[31], i1[31], select);
endmodule